
//`define CORE_TYPE_REDUCED
//`define CORE_TYPE_MINIMAL
//`define CORE_TYPE_CLASSIC_8K
`define CORE_TYPE_CLASSIC_128K
//`define CORE_TYPE_ENCHANCED_8K
//`define CORE_TYPE_ENCHANCED_128K
//`define CORE_TYPE_ENCHANCED_4M
//`define CORE_TYPE_XMEGA


